library IEEE;
use IEEE.std_logic_1164.all;

entity test is 
  
end test;
